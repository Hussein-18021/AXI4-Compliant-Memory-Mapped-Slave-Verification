class Rtransaction;
    


endclass