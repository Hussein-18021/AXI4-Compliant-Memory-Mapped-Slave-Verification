package enuming;
    typedef enum { VALID_BEFORE_READY, READY_BEFORE_VALID } handshake_t;
endpackage