class Rtransaction;

endclass